library ieee;
use ieee.std_logic_1164.all;

package Zifenci_EXT is

    constant FUNCT3_FENCE_I : std_logic_vector(2 downto 0) := b"001";

end package;
