library ieee;
use ieee.std_logic_1164.all;

entity vmem is
end entity;

architecture sim of vmem is
begin



  -- FILE:
  -- addr:data
  --
  --
  --
  --
  p_vmem:
  process
  begin
  end process;

end architecture;
