library ieee;
use ieee.std_logic_1164.all;

package D_EXT is

    constant FUNCT3_D   : std_logic_vector(2 downto 0) := b"011";
    constant FMT2_D     : std_logic_vector(1 downto 0) := b"01";

end package;
