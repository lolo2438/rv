package cnst is

  constant BYTE : natural := 8;

  constant NO_WARNING : boolean := false;

end package;
