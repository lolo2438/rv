package cnst is

  constant BYTE : natural := 8;

end package;
