library ieee;
use ieee.std_logic_1164.all;

entity rv_stb is
end entity;

architecture rtl of rv_stb is
begin
end architecture;
