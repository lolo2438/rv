library ieee;
use ieee.std_logic_1164.all;

package Q_EXT is

    constant FUNCT3_Q        : std_logic_vector(2 downto 0) := b"010";
    constant FMT2_Q          : std_logic_vector(1 downto 0) := b"11";

end package;
